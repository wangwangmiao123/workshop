`timescale 1ns / 1ps

module vga_debug(
	input clk,
	input [31:0] debug_data,
	input [9:0]  h_count,
	input [9:0]  v_count,
	
	output [6:0] debug_addr,
	output [11:0] dout
	
);
	 
endmodule
